LIBRARY ieee ;
USE ieee.stdlogic1164.all ;
ENTITY seg7 IS
	PORT ( bcd    : IN   STDLOGICVECTOR(3 DOWNTO 0) ;\
	leds   : OUT  STDLOGICVECTOR(1 TO 7) ) ;
	END seg7 ;
	
	ARCHITECTURE Behavior OF seg7 IS
	BEGIN
		PROCESS ( bcd )
		BEGIN
			CASE bcd IS      -- abcdefg
			WHEN"0000"   => leds <= "1111110";
			WHEN"0001"   => leds <= "0110000";
			WHEN"0010"   => leds <= "1101101";
			WHEN"0011"   => leds <= "1111001";
			WHEN"0100"   => leds <= "0110011";
			WHEN"0101"   => leds <= "1011011";
			WHEN"0110"   => leds <= "1011111";
			WHEN"0111"   => leds <= "1110000";
			WHEN"1000"   => leds <= "1111111";
			WHEN"1001"   => leds <= "1110011";
			WHEN OTHERS  => leds <= "-------" ;
			END CASE ;
			END PROCESS ;
		END Behavior ;
